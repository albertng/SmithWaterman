`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   15:28:05 06/05/2013
// Design Name:   fifotest
// Module Name:   /afs/cs.stanford.edu/group/evodevo/u/albertng/SmithWaterman/SmithWaterman/firmware/fifotest_tb.v
// Project Name:  m505lx325
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: fifotest
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module fifotest_tb;

	// Inputs
	reg clk;
    reg si_clk;
	reg rst;
	reg [127:0] din;
	reg wr_en;
	reg rd_en;

	// Outputs
	wire [127:0] dout;
	wire full;
	wire empty;

	// Instantiate the Unit Under Test (UUT)
    stream_data_sync_buffer sdsb (
        .rst(rst),
        .wr_clk(si_clk),
        .rd_clk(clk),
        .din(din),
        .wr_en(wr_en),
        .rd_en(rd_en),
        .dout(dout),
        .full(full),
        .empty(empty)
    );

    integer i;
	initial begin
		// Initialize Inputs
		clk = 0;
        si_clk = 0;
		rst = 1;
		din = 0;
		wr_en = 0;
		rd_en = 0;
		#100;
        rst <= 0;
        #100;
        din <= 5;
        wr_en <= 1;
        #10;
        wr_en <= 0;
        #100;
        rd_en <= 1;
        #10;
        rd_en <= 0;
        #100;
        for (i = 0; i < 17; i = i + 1) begin
            wr_en <= 1;
            din <= i + 1;
            #10;
        end
        wr_en <= 0;
        #100;
        for (i = 0; i < 17; i = i + 1) begin
            rd_en <= 1;
            #10;
        end
        rd_en <= 0;
        #200;
        $finish;

	end
    
    always begin
        #5 clk = !clk;
    end
    
    always begin
        #5 si_clk = !si_clk;
    end
    
endmodule

